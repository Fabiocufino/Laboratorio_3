SchemaAssemblaggioCirc1_ottimizzato_unica_terra
C3 0 5 100nF IC=0
R5 1 3 220
R3 4 0 47
R2 4 0 47
C4 0 2 100nF IC=0
R6 3 4 220

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
